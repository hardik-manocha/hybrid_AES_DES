--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:25:15 07/27/2014
-- Design Name:   
-- Module Name:   D:/vlsi/hybrid_aes_des/tb_xor_funct.vhd
-- Project Name:  hybrid_aes_des
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: xor_funct
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_xor_funct IS
END tb_xor_funct;
 
ARCHITECTURE behavior OF tb_xor_funct IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT xor_funct
    PORT(
         a : IN  std_logic_vector(31 downto 0);
         b : IN  std_logic_vector(31 downto 0);
         y : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic_vector(31 downto 0) := (others => '0');
   signal b : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal y : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: xor_funct PORT MAP (
          a => a,
          b => b,
          y => y
        );

   -- Clock process definitions
  -- <clock>_process :process
  -- begin
		--<clock> <= '0';
		---wait for <clock>_period/2;
		--<clock> <= '1';
		--wait for <clock>_period/2;
   --end process;
 

   -- Stimulus process
   process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
				a<="00011010000001101000011010010000";
		wait for 100 ns;
				b<="00110001111111011100010000011100";
     --wait for <clock>_period*10;

      -- insert stimulus here 

     -- wait;
   end process;

END architecture;
